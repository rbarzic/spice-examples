Test ALTERPARAM

.param k1 = 1

V1 1 0 PULSE (0 1 0 100ms 100ms 0 200ms)
R1 1 0 1k
B1 0 3 I=k1*exp(-3*V(1,0))
R3 3 0 1k

.tran 1ms 200ms 1u uic
.options method=gear reltol=1m

.control
   listing e
   run
   alterparam k1=2
   mc_source
   run
   plot tran1.v(3) tran2.v(3) '2000*v(1)'
*   quit
.endc

.end
