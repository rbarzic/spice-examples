* CMOS Inverter testbench for ngspice


.include ./5827_035.lib
.include ./inv_spice.spi




VCC vcc 0 5.0v
*                   TD   TR  TF PW    PER
VX vin 0 pulse 0 5v 20n 10n 10n 100n 200n

.TRAN 10ps 1us

.probe  v(vin) v(vout)
.plot  v(vin) v(vout)

.end

