*******************************
* Begin .SUBCKT model         *
* spice-sdb ver 4.28.2007     *
*******************************
.SUBCKT invx1 A Y vcc gnd 
*==============  Begin SPICE netlist of main design ============
M1 Y A gnd gnd nfet  l=0.18u w=1u
M0 Y A vcc vcc pfet  l=0.18u w=1u
.ends invx1
*******************************
